// first_nios2_system_tb.v

// Generated using ACDS version 12.0 178 at 2013.02.23.21:35:38

`timescale 1 ps / 1 ps
module first_nios2_system_tb (
	);

	wire         first_nios2_system_inst_clk_bfm_clk_clk;                    // first_nios2_system_inst_clk_bfm:clk -> [first_nios2_system_inst:clk_clk, first_nios2_system_inst_reset_bfm:clk]
	wire         first_nios2_system_inst_reset_bfm_reset_reset;              // first_nios2_system_inst_reset_bfm:reset -> first_nios2_system_inst:reset_reset_n
	wire   [9:0] first_nios2_system_inst_led_pio_external_connection_export; // first_nios2_system_inst:led_pio_external_connection_export -> first_nios2_system_inst_led_pio_external_connection_bfm:sig_export
	wire         first_nios2_system_inst_sdram_0_wire_cs_n;                  // first_nios2_system_inst:sdram_0_wire_cs_n -> first_nios2_system_inst_sdram_0_wire_bfm:sig_cs_n
	wire   [1:0] first_nios2_system_inst_sdram_0_wire_ba;                    // first_nios2_system_inst:sdram_0_wire_ba -> first_nios2_system_inst_sdram_0_wire_bfm:sig_ba
	wire   [1:0] first_nios2_system_inst_sdram_0_wire_dqm;                   // first_nios2_system_inst:sdram_0_wire_dqm -> first_nios2_system_inst_sdram_0_wire_bfm:sig_dqm
	wire         first_nios2_system_inst_sdram_0_wire_cke;                   // first_nios2_system_inst:sdram_0_wire_cke -> first_nios2_system_inst_sdram_0_wire_bfm:sig_cke
	wire  [11:0] first_nios2_system_inst_sdram_0_wire_addr;                  // first_nios2_system_inst:sdram_0_wire_addr -> first_nios2_system_inst_sdram_0_wire_bfm:sig_addr
	wire         first_nios2_system_inst_sdram_0_wire_we_n;                  // first_nios2_system_inst:sdram_0_wire_we_n -> first_nios2_system_inst_sdram_0_wire_bfm:sig_we_n
	wire         first_nios2_system_inst_sdram_0_wire_ras_n;                 // first_nios2_system_inst:sdram_0_wire_ras_n -> first_nios2_system_inst_sdram_0_wire_bfm:sig_ras_n
	wire  [15:0] first_nios2_system_inst_sdram_0_wire_dq;                    // [] -> [first_nios2_system_inst:sdram_0_wire_dq, first_nios2_system_inst_sdram_0_wire_bfm:sig_dq]
	wire         first_nios2_system_inst_sdram_0_wire_cas_n;                 // first_nios2_system_inst:sdram_0_wire_cas_n -> first_nios2_system_inst_sdram_0_wire_bfm:sig_cas_n

	first_nios2_system first_nios2_system_inst (
		.clk_clk                            (first_nios2_system_inst_clk_bfm_clk_clk),                    //                         clk.clk
		.reset_reset_n                      (first_nios2_system_inst_reset_bfm_reset_reset),              //                       reset.reset_n
		.led_pio_external_connection_export (first_nios2_system_inst_led_pio_external_connection_export), // led_pio_external_connection.export
		.sdram_0_wire_addr                  (first_nios2_system_inst_sdram_0_wire_addr),                  //                sdram_0_wire.addr
		.sdram_0_wire_ba                    (first_nios2_system_inst_sdram_0_wire_ba),                    //                            .ba
		.sdram_0_wire_cas_n                 (first_nios2_system_inst_sdram_0_wire_cas_n),                 //                            .cas_n
		.sdram_0_wire_cke                   (first_nios2_system_inst_sdram_0_wire_cke),                   //                            .cke
		.sdram_0_wire_cs_n                  (first_nios2_system_inst_sdram_0_wire_cs_n),                  //                            .cs_n
		.sdram_0_wire_dq                    (first_nios2_system_inst_sdram_0_wire_dq),                    //                            .dq
		.sdram_0_wire_dqm                   (first_nios2_system_inst_sdram_0_wire_dqm),                   //                            .dqm
		.sdram_0_wire_ras_n                 (first_nios2_system_inst_sdram_0_wire_ras_n),                 //                            .ras_n
		.sdram_0_wire_we_n                  (first_nios2_system_inst_sdram_0_wire_we_n),                  //                            .we_n
		.sdram_external_clk_clk             ()                                                            //          sdram_external_clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50)
	) first_nios2_system_inst_clk_bfm (
		.clk (first_nios2_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) first_nios2_system_inst_reset_bfm (
		.reset (first_nios2_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (first_nios2_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm first_nios2_system_inst_led_pio_external_connection_bfm (
		.sig_export (first_nios2_system_inst_led_pio_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0002 first_nios2_system_inst_sdram_0_wire_bfm (
		.sig_addr  (first_nios2_system_inst_sdram_0_wire_addr),  // conduit.addr
		.sig_ba    (first_nios2_system_inst_sdram_0_wire_ba),    //        .ba
		.sig_cas_n (first_nios2_system_inst_sdram_0_wire_cas_n), //        .cas_n
		.sig_cke   (first_nios2_system_inst_sdram_0_wire_cke),   //        .cke
		.sig_cs_n  (first_nios2_system_inst_sdram_0_wire_cs_n),  //        .cs_n
		.sig_dq    (first_nios2_system_inst_sdram_0_wire_dq),    //        .dq
		.sig_dqm   (first_nios2_system_inst_sdram_0_wire_dqm),   //        .dqm
		.sig_ras_n (first_nios2_system_inst_sdram_0_wire_ras_n), //        .ras_n
		.sig_we_n  (first_nios2_system_inst_sdram_0_wire_we_n)   //        .we_n
	);

endmodule
