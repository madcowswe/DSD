library verilog;
use verilog.vl_types.all;
entity first_nios2_system_cpu_test_bench is
    port(
        A_bstatus_reg   : in     vl_logic_vector(31 downto 0);
        A_cmp_result    : in     vl_logic;
        A_ctrl_exception: in     vl_logic;
        A_ctrl_ld_non_bypass: in     vl_logic;
        A_dst_regnum    : in     vl_logic_vector(4 downto 0);
        A_en            : in     vl_logic;
        A_estatus_reg   : in     vl_logic_vector(31 downto 0);
        A_ienable_reg   : in     vl_logic_vector(31 downto 0);
        A_ipending_reg  : in     vl_logic_vector(31 downto 0);
        A_iw            : in     vl_logic_vector(31 downto 0);
        A_mem_byte_en   : in     vl_logic_vector(3 downto 0);
        A_op_hbreak     : in     vl_logic;
        A_op_intr       : in     vl_logic;
        A_pcb           : in     vl_logic_vector(24 downto 0);
        A_st_data       : in     vl_logic_vector(31 downto 0);
        A_status_reg    : in     vl_logic_vector(31 downto 0);
        A_valid         : in     vl_logic;
        A_wr_data_unfiltered: in     vl_logic_vector(31 downto 0);
        A_wr_dst_reg    : in     vl_logic;
        E_add_br_to_taken_history_unfiltered: in     vl_logic;
        E_logic_result  : in     vl_logic_vector(31 downto 0);
        E_valid         : in     vl_logic;
        M_bht_ptr_unfiltered: in     vl_logic_vector(7 downto 0);
        M_bht_wr_data_unfiltered: in     vl_logic_vector(1 downto 0);
        M_bht_wr_en_unfiltered: in     vl_logic;
        M_mem_baddr     : in     vl_logic_vector(24 downto 0);
        M_target_pcb    : in     vl_logic_vector(24 downto 0);
        M_valid         : in     vl_logic;
        W_dst_regnum    : in     vl_logic_vector(4 downto 0);
        W_iw            : in     vl_logic_vector(31 downto 0);
        W_iw_op         : in     vl_logic_vector(5 downto 0);
        W_iw_opx        : in     vl_logic_vector(5 downto 0);
        W_pcb           : in     vl_logic_vector(24 downto 0);
        W_valid         : in     vl_logic;
        W_vinst         : in     vl_logic_vector(55 downto 0);
        W_wr_dst_reg    : in     vl_logic;
        clk             : in     vl_logic;
        d_address       : in     vl_logic_vector(24 downto 0);
        d_byteenable    : in     vl_logic_vector(3 downto 0);
        d_read          : in     vl_logic;
        d_write         : in     vl_logic;
        i_address       : in     vl_logic_vector(24 downto 0);
        i_read          : in     vl_logic;
        i_readdatavalid : in     vl_logic;
        reset_n         : in     vl_logic;
        A_wr_data_filtered: out    vl_logic_vector(31 downto 0);
        E_add_br_to_taken_history_filtered: out    vl_logic;
        E_src1_eq_src2  : out    vl_logic;
        M_bht_ptr_filtered: out    vl_logic_vector(7 downto 0);
        M_bht_wr_data_filtered: out    vl_logic_vector(1 downto 0);
        M_bht_wr_en_filtered: out    vl_logic;
        test_has_ended  : out    vl_logic
    );
end first_nios2_system_cpu_test_bench;
