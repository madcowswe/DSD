library verilog;
use verilog.vl_types.all;
entity first_nios2_system_cpu_nios2_performance_monitors is
end first_nios2_system_cpu_nios2_performance_monitors;
