// first_nios2_system_tb.v

// Generated using ACDS version 12.1 177 at 2013.02.26.02:02:36

`timescale 1 ps / 1 ps
module first_nios2_system_tb (
	);

	wire         first_nios2_system_inst_clk_bfm_clk_clk;                    // first_nios2_system_inst_clk_bfm:clk -> [first_nios2_system_inst:clk_clk, first_nios2_system_inst_reset_bfm:clk]
	wire         first_nios2_system_inst_reset_bfm_reset_reset;              // first_nios2_system_inst_reset_bfm:reset -> first_nios2_system_inst:reset_reset_n
	wire   [9:0] first_nios2_system_inst_led_pio_external_connection_export; // first_nios2_system_inst:led_pio_external_connection_export -> first_nios2_system_inst_led_pio_external_connection_bfm:sig_export
	wire         sdram_0_my_partner_clk_bfm_clk_clk;                         // sdram_0_my_partner_clk_bfm:clk -> sdram_0_my_partner:clk
	wire         first_nios2_system_inst_sdram_0_wire_cs_n;                  // first_nios2_system_inst:sdram_0_wire_cs_n -> sdram_0_my_partner:zs_cs_n
	wire   [1:0] first_nios2_system_inst_sdram_0_wire_ba;                    // first_nios2_system_inst:sdram_0_wire_ba -> sdram_0_my_partner:zs_ba
	wire   [1:0] first_nios2_system_inst_sdram_0_wire_dqm;                   // first_nios2_system_inst:sdram_0_wire_dqm -> sdram_0_my_partner:zs_dqm
	wire         first_nios2_system_inst_sdram_0_wire_cke;                   // first_nios2_system_inst:sdram_0_wire_cke -> sdram_0_my_partner:zs_cke
	wire  [11:0] first_nios2_system_inst_sdram_0_wire_addr;                  // first_nios2_system_inst:sdram_0_wire_addr -> sdram_0_my_partner:zs_addr
	wire         first_nios2_system_inst_sdram_0_wire_we_n;                  // first_nios2_system_inst:sdram_0_wire_we_n -> sdram_0_my_partner:zs_we_n
	wire         first_nios2_system_inst_sdram_0_wire_ras_n;                 // first_nios2_system_inst:sdram_0_wire_ras_n -> sdram_0_my_partner:zs_ras_n
	wire         first_nios2_system_inst_sdram_0_wire_cas_n;                 // first_nios2_system_inst:sdram_0_wire_cas_n -> sdram_0_my_partner:zs_cas_n
	wire  [15:0] first_nios2_system_inst_sdram_0_wire_dq;                    // [] -> [first_nios2_system_inst:sdram_0_wire_dq, sdram_0_my_partner:zs_dq]

	first_nios2_system first_nios2_system_inst (
		.clk_clk                            (first_nios2_system_inst_clk_bfm_clk_clk),                    //                         clk.clk
		.reset_reset_n                      (first_nios2_system_inst_reset_bfm_reset_reset),              //                       reset.reset_n
		.led_pio_external_connection_export (first_nios2_system_inst_led_pio_external_connection_export), // led_pio_external_connection.export
		.sdram_0_wire_addr                  (first_nios2_system_inst_sdram_0_wire_addr),                  //                sdram_0_wire.addr
		.sdram_0_wire_ba                    (first_nios2_system_inst_sdram_0_wire_ba),                    //                            .ba
		.sdram_0_wire_cas_n                 (first_nios2_system_inst_sdram_0_wire_cas_n),                 //                            .cas_n
		.sdram_0_wire_cke                   (first_nios2_system_inst_sdram_0_wire_cke),                   //                            .cke
		.sdram_0_wire_cs_n                  (first_nios2_system_inst_sdram_0_wire_cs_n),                  //                            .cs_n
		.sdram_0_wire_dq                    (first_nios2_system_inst_sdram_0_wire_dq),                    //                            .dq
		.sdram_0_wire_dqm                   (first_nios2_system_inst_sdram_0_wire_dqm),                   //                            .dqm
		.sdram_0_wire_ras_n                 (first_nios2_system_inst_sdram_0_wire_ras_n),                 //                            .ras_n
		.sdram_0_wire_we_n                  (first_nios2_system_inst_sdram_0_wire_we_n),                  //                            .we_n
		.clock_bridge_0_out_clk_clk         ()                                                            //      clock_bridge_0_out_clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) first_nios2_system_inst_clk_bfm (
		.clk (first_nios2_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) first_nios2_system_inst_reset_bfm (
		.reset (first_nios2_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (first_nios2_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm first_nios2_system_inst_led_pio_external_connection_bfm (
		.sig_export (first_nios2_system_inst_led_pio_external_connection_export)  // conduit.export
	);

	altera_sdram_partner_module sdram_0_my_partner (
		.clk      (sdram_0_my_partner_clk_bfm_clk_clk),         //     clk.clk
		.zs_dq    (first_nios2_system_inst_sdram_0_wire_dq),    // conduit.dq
		.zs_addr  (first_nios2_system_inst_sdram_0_wire_addr),  //        .addr
		.zs_ba    (first_nios2_system_inst_sdram_0_wire_ba),    //        .ba
		.zs_cas_n (first_nios2_system_inst_sdram_0_wire_cas_n), //        .cas_n
		.zs_cke   (first_nios2_system_inst_sdram_0_wire_cke),   //        .cke
		.zs_cs_n  (first_nios2_system_inst_sdram_0_wire_cs_n),  //        .cs_n
		.zs_dqm   (first_nios2_system_inst_sdram_0_wire_dqm),   //        .dqm
		.zs_ras_n (first_nios2_system_inst_sdram_0_wire_ras_n), //        .ras_n
		.zs_we_n  (first_nios2_system_inst_sdram_0_wire_we_n)   //        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sdram_0_my_partner_clk_bfm (
		.clk (sdram_0_my_partner_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
