// Master custom instruction verilog block
// Instantiates slave altfp modules
// Does add, sub, mul, div
// Interfaces with the nios 2 as an extended (n'd) custom instruction block

/*
altfp_addsub	altfp_addsub_inst (
	.add_sub ( add_sub_sig ),
	.clk_en ( clk_en_sig ),
	.clock ( clock_sig ),
	.dataa ( dataa_sig ),
	.datab ( datab_sig ),
	.result ( result_sig )
	);
*/

//TODO: generate blah

module fp_cust_insn ( 



);

endmodule