library verilog;
use verilog.vl_types.all;
entity altera_merlin_traffic_limiter is
    generic(
        PKT_TRANS_POSTED: integer := 1;
        PKT_DEST_ID_H   : integer := 0;
        PKT_DEST_ID_L   : integer := 0;
        ST_DATA_W       : integer := 72;
        ST_CHANNEL_W    : integer := 32;
        MAX_OUTSTANDING_RESPONSES: integer := 1;
        PIPELINED       : integer := 0;
        ENFORCE_ORDER   : integer := 1;
        PKT_BYTE_CNT_H  : integer := 0;
        PKT_BYTE_CNT_L  : integer := 0;
        PKT_BYTEEN_H    : integer := 0;
        PKT_BYTEEN_L    : integer := 0;
        PKT_TRANS_WRITE : integer := 0;
        PKT_TRANS_READ  : integer := 0;
        VALID_WIDTH     : integer := 1;
        PREVENT_HAZARDS : integer := 0
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        cmd_sink_valid  : in     vl_logic;
        cmd_sink_data   : in     vl_logic_vector;
        cmd_sink_channel: in     vl_logic_vector;
        cmd_sink_startofpacket: in     vl_logic;
        cmd_sink_endofpacket: in     vl_logic;
        cmd_sink_ready  : out    vl_logic;
        cmd_src_valid   : out    vl_logic_vector;
        cmd_src_data    : out    vl_logic_vector;
        cmd_src_channel : out    vl_logic_vector;
        cmd_src_startofpacket: out    vl_logic;
        cmd_src_endofpacket: out    vl_logic;
        cmd_src_ready   : in     vl_logic;
        rsp_sink_valid  : in     vl_logic;
        rsp_sink_data   : in     vl_logic_vector;
        rsp_sink_channel: in     vl_logic_vector;
        rsp_sink_startofpacket: in     vl_logic;
        rsp_sink_endofpacket: in     vl_logic;
        rsp_sink_ready  : out    vl_logic;
        rsp_src_valid   : out    vl_logic;
        rsp_src_data    : out    vl_logic_vector;
        rsp_src_channel : out    vl_logic_vector;
        rsp_src_startofpacket: out    vl_logic;
        rsp_src_endofpacket: out    vl_logic;
        rsp_src_ready   : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PKT_TRANS_POSTED : constant is 1;
    attribute mti_svvh_generic_type of PKT_DEST_ID_H : constant is 1;
    attribute mti_svvh_generic_type of PKT_DEST_ID_L : constant is 1;
    attribute mti_svvh_generic_type of ST_DATA_W : constant is 1;
    attribute mti_svvh_generic_type of ST_CHANNEL_W : constant is 1;
    attribute mti_svvh_generic_type of MAX_OUTSTANDING_RESPONSES : constant is 1;
    attribute mti_svvh_generic_type of PIPELINED : constant is 1;
    attribute mti_svvh_generic_type of ENFORCE_ORDER : constant is 1;
    attribute mti_svvh_generic_type of PKT_BYTE_CNT_H : constant is 1;
    attribute mti_svvh_generic_type of PKT_BYTE_CNT_L : constant is 1;
    attribute mti_svvh_generic_type of PKT_BYTEEN_H : constant is 1;
    attribute mti_svvh_generic_type of PKT_BYTEEN_L : constant is 1;
    attribute mti_svvh_generic_type of PKT_TRANS_WRITE : constant is 1;
    attribute mti_svvh_generic_type of PKT_TRANS_READ : constant is 1;
    attribute mti_svvh_generic_type of VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PREVENT_HAZARDS : constant is 1;
end altera_merlin_traffic_limiter;
