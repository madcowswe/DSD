library verilog;
use verilog.vl_types.all;
entity first_nios2_system_tb is
end first_nios2_system_tb;
